`include "myhead.h"

module csr(
    
);